library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity char_rom is
port (address : in  std_logic_vector(7 downto 0);   -- 256 addresses in total
      data    : out std_logic_vector(63 downto 0));  -- 64 bits/address
end entity;

architecture RTL of char_rom is
begin
process(address)
  begin
  case address is
    --character 1
    when "00000000" => data <= "1111111111111111111111111100000000000000000000000000000000000000";
    when "00000001" => data <= "1111111111111111111111111111111000000000000000000000000000000000";
    when "00000010" => data <= "1111111111111111111111111111111111100000000000000000000000000000";
    when "00000011" => data <= "1111111111111111111111111111111111111110000000000000000000000000";
    when "00000100" => data <= "1111111111110000000000000000011111111111111000000000000000000000";
    when "00000101" => data <= "1111111111110000000000000000011111111111111000000000000000000000";
    when "00000110" => data <= "1111111111110000000000000000011111111111111000000000000000000000";
    when "00000111" => data <= "1111111111110000000000000000011111111111111000000000000000000000";
    when "00001000" => data <= "1111111111110000000000000000011111111111111000000000000000000000";
    when "00001001" => data <= "1111111111110000000000000000011111111111111000000000000000000000";
    when "00001010" => data <= "1111111111110000000000000000011111111111111000000000000000000000";
    when "00001011" => data <= "1111111111110000000000000000011111111111111000000000000000000000";
    when "00001100" => data <= "1111111111110000000000000000011111111111111000000000000000000000";
    when "00001101" => data <= "1111111111110000000000000000011111111111111000000000000000000000";
    when "00001110" => data <= "1111111111110000000000000000011111111111111000000000000000000000";
    when "00001111" => data <= "1111111111110000000000000000011111111111111000000000000000000000";
    when "00010000" => data <= "1111111111110000000000000000011111111111111000000000000000000000";
    when "00010001" => data <= "1111111111110000000000000000011111111111111000000000000000000000";
    when "00010010" => data <= "1111111111110000000000000000011111111111111000000000000000000000";
    when "00010011" => data <= "1111111111110000000000000000011111111111111000000000000000000000";
    when "00010100" => data <= "1111111111110000000000000111111111111110000000000000000000000000";
    when "00010101" => data <= "1111111111110000000001111111111111100000000000000000000000000000";
    when "00010110" => data <= "1111111111110000011111111111111000000000000000000000000000000000";
    when "00010111" => data <= "1111111111111111111111111100000000000000000000000000000000000000";
    when "00011000" => data <= "1111111111111111111111111100000000000000000000000000000000000000";
    when "00011001" => data <= "1111111111111111111111111100000000000000000000000000000000000000";
    when "00011010" => data <= "1111111111111111111111111100000000000000000000000000000000000000";
    when "00011011" => data <= "1111111111111111111111111100000000000000000000000000000000000000";
    when "00011100" => data <= "1111111111110000011111111111111000000000000000000000000000000000";
    when "00011101" => data <= "1111111111110000000001111111111111000000000000000000000000000000";
    when "00011110" => data <= "1111111111110000000001111111111111000000000000000000000000000000";
    when "00011111" => data <= "1111111111110000000000000111111111111000000000000000000000000000";
    when "00100000" => data <= "1111111111110000000000000111111111111100000000000000000000000000";
    when "00100001" => data <= "1111111111110000000000000111111111111110000000000000000000000000";
    when "00100010" => data <= "1111111111110000000000000000011111111111111000000000000000000000";
    when "00100011" => data <= "1111111111110000000000000000000001111111111111100000000000000000";
    when "00100100" => data <= "1111111111110000000000000000000000001111111111111000000000000000";
    when "00100101" => data <= "1111111111110000000000000000000000000001111111111100000000000000";
    when "00100110" => data <= "1111111111110000000000000000000000000001111111111110000000000000";
    when "00100111" => data <= "1111111111110000000000000000000000000001111111111111100000000000";
    when "00101000" => data <= "1111111111110000000000000000000000000000001111111111111000000000";
    when "00101001" => data <= "1111111111110000000000000000000000000000001111111111111100000000";
    when "00101010" => data <= "1111111111110000000000000000000000000000000000111111111111000000";
    when "00101011" => data <= "1111111111110000000000000000000000000000000000111111111111110000";
    when "00101100" => data <= "1111111111110000000000000000000000000000000000001111111111111000";
    when "00101101" => data <= "1111111111110000000000000000000000000000000000001111111111111100";
    when "00101110" => data <= "1111111111110000000000000000000000000000000000000001111111111110";
    when "00101111" => data <= "1111111111110000000000000000000000000000000000000001111111111111";

    --character 2
    when "00110000" => data <= "0000000000001111111111111111111111111111111111111000000000000000";
    when "00110001" => data <= "0000000000001111111111111111111111111111111111111000000000000000";
    when "00110010" => data <= "0000000000001111111111111111111111111111111111111000000000000000";
    when "00110011" => data <= "0000000000001111111111111111111111111111111111111000000000000000";
    when "00110100" => data <= "0000000000001111111111111111111111111111111111111000000000000000";
    when "00110101" => data <= "0000000000001111111111111111111111111111111111111000000000000000";
    when "00110110" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "00110111" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "00111000" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "00111001" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "00111010" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "00111011" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "00111100" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "00111101" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "00111110" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "00111111" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01000000" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01000001" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01000010" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01000011" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01000100" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01000101" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01000110" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01000111" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01001000" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01001001" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01001010" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01001011" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01001100" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01001101" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01001110" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01001111" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01010000" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01010001" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01010010" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01010011" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01010100" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01010101" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01010110" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01010111" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01011000" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01011001" => data <= "0000000000001111111111100000000000000001111111111000000000000000";
    when "01011010" => data <= "0000000000001111111111111111111111111111111111111000000000000000";
    when "01011011" => data <= "0000000000001111111111111111111111111111111111111000000000000000";
    when "01011100" => data <= "0000000000001111111111111111111111111111111111111000000000000000";
    when "01011101" => data <= "0000000000001111111111111111111111111111111111111000000000000000";
    when "01011110" => data <= "0000000000001111111111111111111111111111111111111000000000000000";
    when "01011111" => data <= "0000000000001111111111111111111111111111111111111000000000000000";

    --character 3
    when "01100000" => data <= "1111111111111100000000000000000000000000000000000011111111111111";
    when "01100001" => data <= "1111111111111110000000000000000000000000000000000111111111111111";
    when "01100010" => data <= "1111111111111111000000000000000000000000000000000111111111111111";
    when "01100011" => data <= "1111111111111111100000000000000000000000000000001111111111111111";
    when "01100100" => data <= "1111111111111111110000000000000000000000000000011111111111111111";
    when "01100101" => data <= "1111111111111111111000000000000000000000000000111111111111111111";
    when "01100110" => data <= "1111111111111111111100000000000000000000000001111111111111111111";
    when "01100111" => data <= "1111111111111000111110000000000000000000000111111000111111111111";
    when "01101000" => data <= "1111111111111000011111000000000000000000011111100001111111111111";
    when "01101001" => data <= "1111111111111000011111000000000000000000111111000001111111111111";
    when "01101010" => data <= "1111111111111000011111000000000000000000111111000001111111111111";
    when "01101011" => data <= "1111111111111000011111000000000000000000111111000001111111111111";
    when "01101100" => data <= "1111111111111000011111000000000000000000111111000001111111111111";
    when "01101101" => data <= "1111111111111000011111000000000000000000111111000001111111111111";
    when "01101110" => data <= "1111111111111000011111000000000000000000111111000001111111111111";
    when "01101111" => data <= "1111111111111000011111000000000000000000111111000001111111111111";
    when "01110000" => data <= "1111111111111000011111000000000000000000111111000001111111111111";
    when "01110001" => data <= "1111111111111000011111000000000000000000111111000001111111111111";
    when "01110010" => data <= "1111111111111000011111000000000000000000111111000001111111111111";
    when "01110011" => data <= "1111111111111000011111000000000000000000111111000001111111111111";
    when "01110100" => data <= "1111111111111000011111000000000000000000111111000001111111111111";
    when "01110101" => data <= "1111111111111000001111100000000000000001111110000001111111111111";
    when "01110110" => data <= "1111111111111000000011111000000000000001111100000001111111111111";
    when "01110111" => data <= "1111111111111000000001111100000000000011111000000001111111111111";
    when "01111000" => data <= "1111111111111000000001111100000000000011111000000001111111111111";
    when "01111001" => data <= "1111111111111000000000011111111111111111100000000001111111111111";
    when "01111010" => data <= "1111111111111000000000011111111111111111111000000001111111111111";
    when "01111011" => data <= "1111111111111000000000011111111111111111111000000001111111111111";
    when "01111100" => data <= "1111111111111000000000000000000000000000000000000001111111111111";
    when "01111101" => data <= "1111111111111000000000000000000000000000000000000001111111111111";
    when "01111110" => data <= "1111111111111000000000000000000000000000000000000001111111111111";
    when "01111111" => data <= "1111111111111000000000000000000000000000000000000001111111111111";
    when "10000000" => data <= "1111111111111000000000000000000000000000000000000001111111111111";
    when "10000001" => data <= "1111111111111000000000000000000000000000000000000001111111111111";
    when "10000010" => data <= "1111111111111000000000000000000000000000000000000001111111111111";
    when "10000011" => data <= "1111111111111000000000000000000000000000000000000001111111111111";
    when "10000100" => data <= "1111111111111000000000000000000000000000000000000001111111111111";
    when "10000101" => data <= "1111111111111000000000000000000000000000000000000001111111111111";
    when "10000110" => data <= "1111111111111000000000000000000000000000000000000001111111111111";
    when "10000111" => data <= "1111111111111000000000000000000000000000000000000001111111111111";
    when "10001000" => data <= "1111111111111000000000000000000000000000000000000001111111111111";
    when "10001001" => data <= "1111111111111000000000000000000000000000000000000001111111111111";
    when "10001010" => data <= "1111111111111000000000000000000000000000000000000001111111111111";
    when "10001011" => data <= "1111111111111000000000000000000000000000000000000001111111111111";
    when "10001100" => data <= "1111111111111000000000000000000000000000000000000001111111111111";
    when "10001101" => data <= "1111111111111000000000000000000000000000000000000001111111111111";
    when "10001110" => data <= "1111111111111000000000000000000000000000000000000001111111111111";
    when "10001111" => data <= "1111111111111000000000000000000000000000000000000001111111111111";
    when others => data<= "0000000000000000000000000000000000000000000000000000000000000000";
        -------------------------
 end case;
end process;
end RTL;
